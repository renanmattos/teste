signal a : std_logic;